module util

fn test_auto_id() {
	assert auto_id() > 0
}
