module util

fn test_pair() {
	assert pair(0, ['a', 'b', 'c']).str() == "(0, ['a', 'b', 'c'])"
}
