module util

fn test_tuple() {
	assert tuple2(0, ['a', 'b', 'c']).str() == "(0, ['a', 'b', 'c'])"
}
