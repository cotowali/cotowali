module lsp

// method: ‘textDocument/signatureHelp’
// response: SignatureHelp | none
// request: TextDocumentPositionParams
// struct SymbolInformation {
// }
