// Copyright (c) 2021-2023 zakuro <z@kuro.red>. All rights reserved.
//
// This Source Code Form is subject to the terms of the Mozilla Public
// License, v. 2.0. If a copy of the MPL was not distributed with this
// file, You can obtain one at https://mozilla.org/MPL/2.0/.
module util

fn test_is_relative_path() {
	assert is_relative_path('.')
	assert is_relative_path('./')
	assert is_relative_path('./a')
	assert is_relative_path('../')
	assert is_relative_path('../a')

	assert !is_relative_path('a')
	assert !is_relative_path('/a')
}
