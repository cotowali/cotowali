module sexprs

// TODO

pub struct Emitter {
	builder code.Builder
}
