// Copyright (c) 2021 zakuro <z@kuro.red>. All rights reserved.
//
// This Source Code Form is subject to the terms of the Mozilla Public
// License, v. 2.0. If a copy of the MPL was not distributed with this
// file, You can obtain one at https://mozilla.org/MPL/2.0/.
module symbols

import cotowali.errors { unreachable }

pub struct RegisterFnArgs {
	Var
	FunctionTypeInfo
}

pub struct FunctionTypeInfo {
pub:
	receiver Type = builtin_type(.placeholder)
	pipe_in  Type = builtin_type(.void)
	params   []Type
	ret      Type = builtin_type(.void)
}

pub fn (ts TypeSymbol) function_info() ?FunctionTypeInfo {
	resolved := ts.resolved()
	return if resolved.info is FunctionTypeInfo { resolved.info } else { none }
}

pub fn (f &FunctionTypeInfo) is_method() bool {
	return f.receiver != builtin_type(.placeholder)
}

fn (f &FunctionTypeInfo) signature(s &Scope) string {
	params_str := f.params.map(s.must_lookup_type(it).name).join(', ')
	in_str := s.must_lookup_type(f.pipe_in).name
	ret_str := s.must_lookup_type(f.ret).name

	return (if f.is_method() {
		'fn (${s.must_lookup_type(f.receiver).name})'
	} else {
		'fn'
	}) + ' $in_str | ($params_str) $ret_str'
}

pub fn (t TypeSymbol) fn_signature() ?string {
	return if t.info is FunctionTypeInfo {
		t.info.signature(t.scope() or { panic(unreachable(err)) })
	} else {
		none
	}
}

pub fn (mut s Scope) lookup_or_register_fn_type(info FunctionTypeInfo) &TypeSymbol {
	typename := info.signature(s)
	return s.lookup_or_register_type(name: typename, info: info)
}

pub fn (s Scope) lookup_fn_type(info FunctionTypeInfo) ?&TypeSymbol {
	typename := info.signature(s)
	return s.lookup_type(typename)
}

pub fn (mut s Scope) register_fn(f RegisterFnArgs) ?&Var {
	typ := s.lookup_or_register_fn_type(f.FunctionTypeInfo).typ
	return s.register_var(Var{ ...f.Var, typ: typ })
}

fn (mut s Scope) must_register_fn(f RegisterFnArgs) &Var {
	return s.register_fn(f) or { panic(unreachable(err)) }
}

// -- methods --

pub fn (mut s Scope) register_method(f RegisterFnArgs) ?&Var {
	if !f.is_method() {
		panic(unreachable('not a method'))
	}
	typ := s.lookup_or_register_fn_type(f.FunctionTypeInfo).typ
	v := &Var{
		...f.Var
		id: if f.Var.id == 0 { auto_id() } else { f.Var.id }
		typ: typ
		receiver_typ: f.FunctionTypeInfo.receiver
		scope: s
	}
	if v.name in s.methods[typ] {
		return error('duplicated method $v.name')
	}
	s.methods[typ][v.name] = s
	return v
}

pub fn (mut s Scope) lookup_method(typ Type, name string) ?&Var {
	return (s.methods[typ] or { return none })[name] or { return none }
}
