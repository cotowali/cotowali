// Copyright (c) 2021 The Cotowali Authors. All rights reserved.
//
// This Source Code Form is subject to the terms of the Mozilla Public
// License, v. 2.0. If a copy of the MPL was not distributed with this
// file, You can obtain one at https://mozilla.org/MPL/2.0/.
module sh

import cotowali.ast { MapLiteral }

fn (mut e Emitter) map_literal(expr MapLiteral, opt ExprOpt) {
	panic('unimplemented')
}
