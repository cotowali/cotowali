module types

struct TypeSymbol {
pub:
	name string
}
