module emit

import cotowari.ast { Pipeline, Stmt }
import cotowari.symbols

pub fn (mut g Gen) gen(f ast.File) {
	g.file(f)
}

fn (mut g Gen) file(f ast.File) {
	g.builtin()
	g.writeln('# file: $f.path')
	g.stmts(f.stmts)
}

fn (mut g Gen) builtin() {
	f := $embed_file('../../builtin/builtin.sh')
	g.writeln(f.to_string())
}

fn (mut g Gen) stmts(stmts []Stmt) {
	for stmt in stmts {
		g.stmt(stmt)
	}
}

fn (mut g Gen) stmt(stmt Stmt) {
	match stmt {
		ast.FnDecl {
			g.fn_decl(stmt)
		}
		ast.Block {
			g.block(stmt)
		}
		ast.Expr {
			g.expr(stmt, as_command: true, writeln: true)
		}
		ast.AssignStmt {
			g.assign(stmt)
		}
		ast.EmptyStmt {
			g.writeln('')
		}
		ast.ForInStmt {
			g.for_in_stmt(stmt)
		}
		ast.IfStmt {
			g.if_stmt(stmt)
		}
	}
}

fn (mut g Gen) block(block ast.Block) {
	g.stmts(block.stmts)
}

fn (mut g Gen) if_stmt(stmt ast.IfStmt) {
	for i, branch in stmt.branches {
		mut is_else := i == stmt.branches.len - 1 && stmt.has_else
		if is_else {
			g.writeln('else')
		} else {
			g.write(if i == 0 { 'if ' } else { 'elif ' })
			g.expr(branch.cond, as_command: true, writeln: true)
			g.writeln('then')
		}
		g.indent++
		g.block(branch.body)
		g.indent--
	}
	g.writeln('fi')
}

fn (mut g Gen) for_in_stmt(stmt ast.ForInStmt) {
	g.write('for $stmt.val.full_name() in ')
	g.expr(stmt.expr, writeln: true)
	g.writeln('do')
	g.indent++
	g.block(stmt.body)
	g.indent--
	g.writeln('done')
}

struct ExprOpt {
	as_command bool
	writeln    bool
}

fn (mut g Gen) expr(expr ast.Expr, opt ExprOpt) {
	match expr {
		ast.CallFn {
			g.call_fn(expr, opt)
		}
		ast.Pipeline {
			g.pipeline(expr, opt)
		}
		ast.InfixExpr {
			g.infix_expr(expr, opt)
		}
		ast.IntLiteral {
			if opt.as_command {
				g.write('echo ')
			}
			g.write(expr.token.text)
		}
		symbols.Var {
			if opt.as_command {
				g.write('echo ')
			}
			g.write('"\$$expr.full_name()"')
		}
	}
	if opt.writeln {
		g.writeln('')
	}
}

fn (mut g Gen) infix_expr(expr ast.InfixExpr, opt ExprOpt) {
	op := expr.op
	match op.kind {
		.op_plus, .op_minus, .op_div, .op_mul {
			if opt.as_command {
				g.write('echo ')
			}
			g.write('\$(( (')
			g.expr(expr.left, {})
			g.write(' $op.text ')
			g.expr(expr.right, {})
			g.write(') ))')
		}
		else {
			panic('unimplemented')
		}
	}
}

fn (mut g Gen) pipeline(stmt Pipeline, opt ExprOpt) {
	if !opt.as_command {
		g.write('\$(')
	}

	for i, expr in stmt.exprs {
		if i > 0 {
			g.write(' | ')
		}
		g.expr(expr, as_command: true)
	}
	g.writeln('')

	if !opt.as_command {
		g.write(')')
	}
}

fn (mut g Gen) call_fn(expr ast.CallFn, opt ExprOpt) {
	if !opt.as_command {
		g.write('\$(')
	}

	g.write(expr.func.full_name())
	for arg in expr.args {
		g.write(' ')
		g.expr(arg, {})
	}

	if !opt.as_command {
		g.write(')')
	}
}

fn (mut g Gen) fn_decl(node ast.FnDecl) {
	g.writeln('${node.name}() {')
	g.indent++
	for i, param in node.params {
		g.writeln('$param.full_name()=\$${i + 1}')
	}
	g.block(node.body)
	g.indent--
	g.writeln('}')
}

fn (mut g Gen) assign(node ast.AssignStmt) {
	g.write('$node.left.full_name()=')
	g.expr(node.right, {})
	g.writeln('')
}
