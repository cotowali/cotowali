module checker

import cotowari.ast

pub fn (c Checker) check_file(mut f ast.File) {
}
