module ast

pub struct File {
pub:
	path string
}
