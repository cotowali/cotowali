module lsp

// method: ‘textDocument/implementation’
// response: Location | []Location | []LocationLink | none
// request: TextDocumentPositionParams
