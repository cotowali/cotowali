module config

[heap]
pub struct Config {
}

pub fn new_config() &Config {
	return {}
}
